module c

#flag -I @VMODROOT/HieroglyphVM/src
#include "chunk.h"
